`ifndef DEFINE
`define DEFINE

parameter XLEN = 32;

parameter PC_START_ADDR = 32'h00000000;
parameter SP_START_ADDR = 32'h0000FFFE;

parameter IMEM_SIZE = 65536; // 64 KB
parameter DMEM_SIZE = 65536; // 64 KB

`endif
