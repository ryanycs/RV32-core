module mul (
    input  logic  clk,
    input  logic  rst,

    input  logic [31:0]  a,
    input  logic [31:0]  b,
    input  logic         mul_ctrl,
    output logic [63:0]  mul_result
);

endmodule
